`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.06.2025 19:37:17
// Design Name: 
// Module Name: set_associative_fifo
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module set_associative_fifo(
  input clk, reset,
  input cpu_req, cpu_write,
  input [31:0] cpu_addr,
  input [31:0] cpu_write_data,
  output reg [31:0] cpu_read_data,
  output reg hit1, hit2, hit3, hit4,
  output reg HIT, MISS,
  output reg mem_req, mem_write,
  output reg [31:0] mem_addr,
  output reg [31:0] mem_write_data,
  input [31:0] mem_read_data,
  // --- ADDED THESE OUTPUT PORTS ---
  output reg [1:0] fifo_counter_out,
  output reg [31:0] hit_count,
  output reg [31:0] miss_count
);

  reg [255:0] valid1, valid2, valid3, valid4;
  reg [21:0] tag1[0:255], tag2[0:255], tag3[0:255], tag4[0:255];
  reg [31:0] data1[0:255], data2[0:255], data3[0:255], data4[0:255];
  reg [1:0] fifo_counter[0:255];

  // Combinational signals based on current cpu_addr
  wire [21:0] tag = cpu_addr[31:10];
  wire [7:0] index = cpu_addr[9:2];

  // Combinational hit checks for each way
  wire cache_hit1_comb = (valid1[index] == 1'b1) && (tag1[index] == tag);
  wire cache_hit2_comb = (valid2[index] == 1'b1) && (tag2[index] == tag);
  wire cache_hit3_comb = (valid3[index] == 1'b1) && (tag3[index] == tag);
  wire cache_hit4_comb = (valid4[index] == 1'b1) && (tag4[index] == tag);

  // Overall combinatorial hit
  wire cache_hit_comb = cache_hit1_comb || cache_hit2_comb || cache_hit3_comb || cache_hit4_comb;

  // Registered internal values for outputs
  reg [31:0] hit_count_internal; // Renamed to avoid clash with port name
  reg [31:0] miss_count_internal; // Renamed
  reg [1:0] fifo_counter_out_internal; // Renamed

  // Output assignments to reflect internal registered values
  // Since the output ports are now declared as 'reg', we directly assign to them.
  // The 'assign' statement would be for 'wire' outputs.
  // We'll directly assign to the output regs inside the always block.


  integer i;

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      for(i = 0; i < 256; i = i + 1) begin
        valid1[i] <= 0; valid2[i] <= 0; valid3[i] <= 0; valid4[i] <= 0;
        tag1[i] <= 0; tag2[i] <= 0; tag3[i] <= 0; tag4[i] <= 0;
        data1[i] <= 0; data2[i] <= 0; data3[i] <= 0; data4[i] <= 0;
        fifo_counter[i] <= 0;
      end
      hit1 <= 0; hit2 <= 0; hit3 <= 0; hit4 <= 0; HIT <= 0; MISS <= 0;
      mem_req <= 0; mem_write <= 0;
      mem_addr <= 0; mem_write_data <= 0;
      cpu_read_data <= 0;
      hit_count <= 0; // Directly assign to output reg
      miss_count <= 0; // Directly assign to output reg
      fifo_counter_out <= 0; // Directly assign to output reg
    end
    else begin
      // Default de-assertion for single-cycle control signals
      mem_req <= 0;
      mem_write <= 0;
      HIT <= 0;
      MISS <= 0;
      hit1 <= 0; hit2 <= 0; hit3 <= 0; hit4 <= 0;
      cpu_read_data <= 0; // Clear read data by default unless assigned below

      if(cpu_req) begin
        hit1 <= cache_hit1_comb;
        hit2 <= cache_hit2_comb;
        hit3 <= cache_hit3_comb;
        hit4 <= cache_hit4_comb;
        HIT <= cache_hit_comb;
        MISS <= ~cache_hit_comb;

        if(cache_hit_comb) begin
          hit_count <= hit_count + 1; // Direct update to output reg

          if(!cpu_write) begin // Read hit
            if(cache_hit1_comb) cpu_read_data <= data1[index];
            else if(cache_hit2_comb) cpu_read_data <= data2[index];
            else if(cache_hit3_comb) cpu_read_data <= data3[index];
            else if(cache_hit4_comb) cpu_read_data <= data4[index];
          end else begin // Write hit
            mem_req <= 1; // Write-through cache
            mem_write <= 1;
            mem_addr <= cpu_addr;
            mem_write_data <= cpu_write_data;

            if(cache_hit1_comb) data1[index] <= cpu_write_data;
            else if(cache_hit2_comb) data2[index] <= cpu_write_data;
            else if(cache_hit3_comb) data3[index] <= cpu_write_data;
            else if(cache_hit4_comb) data4[index] <= cpu_write_data;
          end
        end else begin // Miss
          miss_count <= miss_count + 1; // Direct update to output reg
          mem_req <= 1;
          mem_addr <= cpu_addr;

          if(cpu_write) begin // Write miss
            mem_write <= 1;
            mem_write_data <= cpu_write_data;
            case(fifo_counter[index])
              2'd0: begin data1[index] <= cpu_write_data; tag1[index] <= tag; valid1[index] <= 1; end
              2'd1: begin data2[index] <= cpu_write_data; tag2[index] <= tag; valid2[index] <= 1; end
              2'd2: begin data3[index] <= cpu_write_data; tag3[index] <= tag; valid3[index] <= 1; end
              2'd3: begin data4[index] <= cpu_write_data; tag4[index] <= tag; valid4[index] <= 1; end
            endcase
          end else begin // Read miss
            cpu_read_data <= mem_read_data; // This means mem_read_data must be valid in the same cycle
            case(fifo_counter[index])
              2'd0: begin data1[index] <= mem_read_data; tag1[index] <= tag; valid1[index] <= 1; end
              2'd1: begin data2[index] <= mem_read_data; tag2[index] <= tag; valid2[index] <= 1; end
              2'd2: begin data3[index] <= mem_read_data; tag3[index] <= tag; valid3[index] <= 1; end
              2'd3: begin data4[index] <= mem_read_data; tag4[index] <= tag; valid4[index] <= 1; end
            endcase
          end
          fifo_counter[index] <= (fifo_counter[index] == 3) ? 0 : fifo_counter[index] + 1;
        end
      end
      // Update fifo_counter_out based on the index currently being processed
      fifo_counter_out <= fifo_counter[index]; // Direct update to output reg
    end
  end
endmodule